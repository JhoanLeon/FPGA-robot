/*
Created by: Jhoan Esteban Leon - je.leon.e@outlook.com
with libraries from https://github.com/freecores/verilog_fixed_point_math_library

inputs and output are in fixed point 17b notation U(17,8) U(N,Q)
*/

//=======================================================
//  MODULE Definition
//=======================================================

module POS_CONTROLLER
(
	//////////// INPUTS //////////
	POS_CONTROLLER_TARGETX_InBus,
	POS_CONTROLLER_TARGETY_InBus,
	POS_CONTROLLER_TARGETTHETA_InBus,
	
	POS_CONTROLLER_CURRENTX_InBus,
	POS_CONTROLLER_CURRENTY_InBus,
	POS_CONTROLLER_CURRENTTHETA_InBus,
	
	//////////// OUTPUTS //////////
	POS_CONTROLLER_GOAL_OutLow, // flag to indicate that the goal is reached
	
	POS_CONTROLLER_ERROR_X_OutBus,
	POS_CONTROLLER_ERROR_Y_OutBus,
	
	POS_CONTROLLER_VX_OutBus,
	POS_CONTROLLER_VY_OutBus,
	POS_CONTROLLER_WZ_OutBus
);

//=======================================================
//  PARAMETER declarations
//=======================================================
parameter N_WIDTH = 17;
parameter Q_WIDTH = 8;

//=======================================================
//  PORT declarations
//=======================================================
input [N_WIDTH-1:0]	POS_CONTROLLER_TARGETX_InBus;
input [N_WIDTH-1:0]	POS_CONTROLLER_TARGETY_InBus;
input [N_WIDTH-1:0]	POS_CONTROLLER_TARGETTHETA_InBus;
	
input [N_WIDTH-1:0]	POS_CONTROLLER_CURRENTX_InBus;
input [N_WIDTH-1:0]	POS_CONTROLLER_CURRENTY_InBus;
input [N_WIDTH-1:0]	POS_CONTROLLER_CURRENTTHETA_InBus;

output POS_CONTROLLER_GOAL_OutLow;

output [N_WIDTH-1:0]	POS_CONTROLLER_ERROR_X_OutBus;
output [N_WIDTH-1:0]	POS_CONTROLLER_ERROR_Y_OutBus;
	
output [N_WIDTH-1:0]	POS_CONTROLLER_VX_OutBus;
output [N_WIDTH-1:0]	POS_CONTROLLER_VY_OutBus;
output [N_WIDTH-1:0]	POS_CONTROLLER_WZ_OutBus;

//=======================================================
//  REG/WIRE declarations
//=======================================================
wire [N_WIDTH-1:0] error_pos_x;
wire [N_WIDTH-1:0] error_pos_y;
wire [N_WIDTH-1:0] error_theta;

//=======================================================
//  STRUCTURAL coding
//=======================================================

qadd #(.Q(Q_WIDTH), .N(N_WIDTH)) sub_error_x
(
    .a(POS_CONTROLLER_TARGETX_InBus),
    .b({~POS_CONTROLLER_CURRENTX_InBus[N_WIDTH-1],POS_CONTROLLER_CURRENTX_InBus[N_WIDTH-2:0]}),
    .c(error_pos_x)
);


qadd #(.Q(Q_WIDTH), .N(N_WIDTH)) sub_error_y
(
    .a(POS_CONTROLLER_TARGETY_InBus),
    .b({~POS_CONTROLLER_CURRENTY_InBus[N_WIDTH-1],POS_CONTROLLER_CURRENTY_InBus[N_WIDTH-2:0]}),
    .c(error_pos_y)
);


qadd #(.Q(Q_WIDTH), .N(N_WIDTH)) sub_error_theta
(
    .a(POS_CONTROLLER_TARGETTHETA_InBus),
    .b({~POS_CONTROLLER_CURRENTTHETA_InBus[N_WIDTH-1],POS_CONTROLLER_CURRENTTHETA_InBus[N_WIDTH-2:0]}),
    .c(error_theta)
);


ERROR_CONTROL error_management
(
	//////////// INPUTS //////////
	.ERROR_CONTROL_X_InBus(error_pos_x),
	.ERROR_CONTROL_Y_InBus(error_pos_y),
	.ERROR_CONTROL_Z_InBus(error_theta),
	
	//////////// OUTPUTS //////////
	.ERROR_CONTROL_GOAL_FLAG(POS_CONTROLLER_GOAL_OutLow),
	
	.ERROR_CONTROL_VX_OutBus(POS_CONTROLLER_VX_OutBus), 
	.ERROR_CONTROL_VY_OutBus(POS_CONTROLLER_VY_OutBus), 
	.ERROR_CONTROL_WZ_OutBus(POS_CONTROLLER_WZ_OutBus) 
);


assign POS_CONTROLLER_ERROR_X_OutBus = error_pos_x;
assign POS_CONTROLLER_ERROR_Y_OutBus = error_pos_y;

endmodule
